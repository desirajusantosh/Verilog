module test();
